module Filter_161Tap(
	input clk,
	//input [19:0]in,
	input [39:0]in,
	input [15:0] h0,
	input [15:0] h1,
	input [15:0] h2,
	input [15:0] h3,
	input [15:0] h4,
	input [15:0] h5,
	input [15:0] h6,
	input [15:0] h7,
	input [15:0] h8,
	input [15:0] h9,
	input [15:0] h10,
	input [15:0] h11,
	input [15:0] h12,
	input [15:0] h13,
	input [15:0] h14,
	input [15:0] h15,
	input [15:0] h16,
	input [15:0] h17,
	input [15:0] h18,
	input [15:0] h19,
	input [15:0] h20,
	input [15:0] h21,
	input [15:0] h22,
	input [15:0] h23,
	input [15:0] h24,
	input [15:0] h25,
	input [15:0] h26,
	input [15:0] h27,
	input [15:0] h28,
	input [15:0] h29,
	input [15:0] h30,
	input [15:0] h31,
	input [15:0] h32,
	input [15:0] h33,
	input [15:0] h34,
	input [15:0] h35,
	input [15:0] h36,
	input [15:0] h37,
	input [15:0] h38,
	input [15:0] h39,
	input [15:0] h40,
	input [15:0] h41,
	input [15:0] h42,
	input [15:0] h43,
	input [15:0] h44,
	input [15:0] h45,
	input [15:0] h46,
	input [15:0] h47,
	input [15:0] h48,
	input [15:0] h49,
	input [15:0] h50,
	input [15:0] h51,
	input [15:0] h52,
	input [15:0] h53,
	input [15:0] h54,
	input [15:0] h55,
	input [15:0] h56,
	input [15:0] h57,
	input [15:0] h58,
	input [15:0] h59,
	input [15:0] h60,
	input [15:0] h61,
	input [15:0] h62,
	input [15:0] h63,
	input [15:0] h64,
	input [15:0] h65,
	input [15:0] h66,
	input [15:0] h67,
	input [15:0] h68,
	input [15:0] h69,
	input [15:0] h70,
	input [15:0] h71,
	input [15:0] h72,
	input [15:0] h73,
	input [15:0] h74,
	input [15:0] h75,
	input [15:0] h76,
	input [15:0] h77,
	input [15:0] h78,
	input [15:0] h79,
	input [15:0] h80,
	output [39:0] out
);

wire [19:0] z0;
wire [19:0] z1;
wire [19:0] z2;
wire [19:0] z3;
wire [19:0] z4;
wire [19:0] z5;
wire [19:0] z6;
wire [19:0] z7;
wire [19:0] z8;
wire [19:0] z9;
wire [19:0] z10;
wire [19:0] z11;
wire [19:0] z12;
wire [19:0] z13;
wire [19:0] z14;
wire [19:0] z15;
wire [19:0] z16;
wire [19:0] z17;
wire [19:0] z18;
wire [19:0] z19;
wire [19:0] z20;
wire [19:0] z21;
wire [19:0] z22;
wire [19:0] z23;
wire [19:0] z24;
wire [19:0] z25;
wire [19:0] z26;
wire [19:0] z27;
wire [19:0] z28;
wire [19:0] z29;
wire [19:0] z30;
wire [19:0] z31;
wire [19:0] z32;
wire [19:0] z33;
wire [19:0] z34;
wire [19:0] z35;
wire [19:0] z36;
wire [19:0] z37;
wire [19:0] z38;
wire [19:0] z39;
wire [19:0] z40;
wire [19:0] z41;
wire [19:0] z42;
wire [19:0] z43;
wire [19:0] z44;
wire [19:0] z45;
wire [19:0] z46;
wire [19:0] z47;
wire [19:0] z48;
wire [19:0] z49;
wire [19:0] z50;
wire [19:0] z51;
wire [19:0] z52;
wire [19:0] z53;
wire [19:0] z54;
wire [19:0] z55;
wire [19:0] z56;
wire [19:0] z57;
wire [19:0] z58;
wire [19:0] z59;
wire [19:0] z60;
wire [19:0] z61;
wire [19:0] z62;
wire [19:0] z63;
wire [19:0] z64;
wire [19:0] z65;
wire [19:0] z66;
wire [19:0] z67;
wire [19:0] z68;
wire [19:0] z69;
wire [19:0] z70;
wire [19:0] z71;
wire [19:0] z72;
wire [19:0] z73;
wire [19:0] z74;
wire [19:0] z75;
wire [19:0] z76;
wire [19:0] z77;
wire [19:0] z78;
wire [19:0] z79;
wire [19:0] z80;
wire [19:0] z81;
wire [19:0] z82;
wire [19:0] z83;
wire [19:0] z84;
wire [19:0] z85;
wire [19:0] z86;
wire [19:0] z87;
wire [19:0] z88;
wire [19:0] z89;
wire [19:0] z90;
wire [19:0] z91;
wire [19:0] z92;
wire [19:0] z93;
wire [19:0] z94;
wire [19:0] z95;
wire [19:0] z96;
wire [19:0] z97;
wire [19:0] z98;
wire [19:0] z99;
wire [19:0] z100;
wire [19:0] z101;
wire [19:0] z102;
wire [19:0] z103;
wire [19:0] z104;
wire [19:0] z105;
wire [19:0] z106;
wire [19:0] z107;
wire [19:0] z108;
wire [19:0] z109;
wire [19:0] z110;
wire [19:0] z111;
wire [19:0] z112;
wire [19:0] z113;
wire [19:0] z114;
wire [19:0] z115;
wire [19:0] z116;
wire [19:0] z117;
wire [19:0] z118;
wire [19:0] z119;
wire [19:0] z120;
wire [19:0] z121;
wire [19:0] z122;
wire [19:0] z123;
wire [19:0] z124;
wire [19:0] z125;
wire [19:0] z126;
wire [19:0] z127;
wire [19:0] z128;
wire [19:0] z129;
wire [19:0] z130;
wire [19:0] z131;
wire [19:0] z132;
wire [19:0] z133;
wire [19:0] z134;
wire [19:0] z135;
wire [19:0] z136;
wire [19:0] z137;
wire [19:0] z138;
wire [19:0] z139;
wire [19:0] z140;
wire [19:0] z141;
wire [19:0] z142;
wire [19:0] z143;
wire [19:0] z144;
wire [19:0] z145;
wire [19:0] z146;
wire [19:0] z147;
wire [19:0] z148;
wire [19:0] z149;
wire [19:0] z150;
wire [19:0] z151;
wire [19:0] z152;
wire [19:0] z153;
wire [19:0] z154;
wire [19:0] z155;
wire [19:0] z156;
wire [19:0] z157;
wire [19:0] z158;
wire [19:0] z159;
wire [19:0] z160;

reg [29:0] add0;
reg [29:0] add1;
reg [29:0] add2;
reg [29:0] add3;
reg [29:0] add4;
reg [29:0] add5;
reg [29:0] add6;
reg [29:0] add7;
reg [29:0] add8;
reg [29:0] add9;
reg [29:0] add10;
reg [29:0] add11;
reg [29:0] add12;
reg [29:0] add13;
reg [29:0] add14;
reg [29:0] add15;
reg [29:0] add16;
reg [29:0] add17;
reg [29:0] add18;
reg [29:0] add19;
reg [29:0] add20;
reg [29:0] add21;
reg [29:0] add22;
reg [29:0] add23;
reg [29:0] add24;
reg [29:0] add25;
reg [29:0] add26;
reg [29:0] add27;
reg [29:0] add28;
reg [29:0] add29;
reg [29:0] add30;
reg [29:0] add31;
reg [29:0] add32;
reg [29:0] add33;
reg [29:0] add34;
reg [29:0] add35;
reg [29:0] add36;
reg [29:0] add37;
reg [29:0] add38;
reg [29:0] add39;
reg [29:0] add40;
reg [29:0] add41;
reg [29:0] add42;
reg [29:0] add43;
reg [29:0] add44;
reg [29:0] add45;
reg [29:0] add46;
reg [29:0] add47;
reg [29:0] add48;
reg [29:0] add49;
reg [29:0] add50;
reg [29:0] add51;
reg [29:0] add52;
reg [29:0] add53;
reg [29:0] add54;
reg [29:0] add55;
reg [29:0] add56;
reg [29:0] add57;
reg [29:0] add58;
reg [29:0] add59;
reg [29:0] add60;
reg [29:0] add61;
reg [29:0] add62;
reg [29:0] add63;
reg [29:0] add64;
reg [29:0] add65;
reg [29:0] add66;
reg [29:0] add67;
reg [29:0] add68;
reg [29:0] add69;
reg [29:0] add70;
reg [29:0] add71;
reg [29:0] add72;
reg [29:0] add73;
reg [29:0] add74;
reg [29:0] add75;
reg [29:0] add76;
reg [29:0] add77;
reg [29:0] add78;
reg [29:0] add79;

reg [39:0] mult0;
reg [39:0] mult1;
reg [39:0] mult2;
reg [39:0] mult3;
reg [39:0] mult4;
reg [39:0] mult5;
reg [39:0] mult6;
reg [39:0] mult7;
reg [39:0] mult8;
reg [39:0] mult9;
reg [39:0] mult10;
reg [39:0] mult11;
reg [39:0] mult12;
reg [39:0] mult13;
reg [39:0] mult14;
reg [39:0] mult15;
reg [39:0] mult16;
reg [39:0] mult17;
reg [39:0] mult18;
reg [39:0] mult19;
reg [39:0] mult20;
reg [39:0] mult21;
reg [39:0] mult22;
reg [39:0] mult23;
reg [39:0] mult24;
reg [39:0] mult25;
reg [39:0] mult26;
reg [39:0] mult27;
reg [39:0] mult28;
reg [39:0] mult29;
reg [39:0] mult30;
reg [39:0] mult31;
reg [39:0] mult32;
reg [39:0] mult33;
reg [39:0] mult34;
reg [39:0] mult35;
reg [39:0] mult36;
reg [39:0] mult37;
reg [39:0] mult38;
reg [39:0] mult39;
reg [39:0] mult40;
reg [39:0] mult41;
reg [39:0] mult42;
reg [39:0] mult43;
reg [39:0] mult44;
reg [39:0] mult45;
reg [39:0] mult46;
reg [39:0] mult47;
reg [39:0] mult48;
reg [39:0] mult49;
reg [39:0] mult50;
reg [39:0] mult51;
reg [39:0] mult52;
reg [39:0] mult53;
reg [39:0] mult54;
reg [39:0] mult55;
reg [39:0] mult56;
reg [39:0] mult57;
reg [39:0] mult58;
reg [39:0] mult59;
reg [39:0] mult60;
reg [39:0] mult61;
reg [39:0] mult62;
reg [39:0] mult63;
reg [39:0] mult64;
reg [39:0] mult65;
reg [39:0] mult66;
reg [39:0] mult67;
reg [39:0] mult68;
reg [39:0] mult69;
reg [39:0] mult70;
reg [39:0] mult71;
reg [39:0] mult72;
reg [39:0] mult73;
reg [39:0] mult74;
reg [39:0] mult75;
reg [39:0] mult76;
reg [39:0] mult77;
reg [39:0] mult78;
reg [39:0] mult79;
reg [39:0] mult80;

reg [39:0] add_0;
reg [39:0] add_1;
reg [39:0] add_2;
reg [39:0] add_3;
reg [39:0] add_4;
reg [39:0] add_5;
reg [39:0] add_6;
reg [39:0] add_7;
reg [39:0] add_8;
reg [39:0] add_9;
reg [39:0] add_10;
reg [39:0] add_11;
reg [39:0] add_12;
reg [39:0] add_13;
reg [39:0] add_14;
reg [39:0] add_15;
reg [39:0] add_16;
reg [39:0] add_17;
reg [39:0] add_18;
reg [39:0] add_19;
reg [39:0] add_20;
reg [39:0] add_21;
reg [39:0] add_22;
reg [39:0] add_23;
reg [39:0] add_24;
reg [39:0] add_25;
reg [39:0] add_26;
reg [39:0] add_27;
reg [39:0] add_28;
reg [39:0] add_29;
reg [39:0] add_30;
reg [39:0] add_31;
reg [39:0] add_32;
reg [39:0] add_33;
reg [39:0] add_34;
reg [39:0] add_35;
reg [39:0] add_36;
reg [39:0] add_37;
reg [39:0] add_38;
reg [39:0] add_39;
reg [39:0] add_40;
reg [39:0] add_41;
reg [39:0] add_42;
reg [39:0] add_43;
reg [39:0] add_44;
reg [39:0] add_45;
reg [39:0] add_46;
reg [39:0] add_47;
reg [39:0] add_48;
reg [39:0] add_49;
reg [39:0] add_50;
reg [39:0] add_51;
reg [39:0] add_52;
reg [39:0] add_53;
reg [39:0] add_54;
reg [39:0] add_55;
reg [39:0] add_56;
reg [39:0] add_57;
reg [39:0] add_58;
reg [39:0] add_59;
reg [39:0] add_60;
reg [39:0] add_61;
reg [39:0] add_62;
reg [39:0] add_63;
reg [39:0] add_64;
reg [39:0] add_65;
reg [39:0] add_66;
reg [39:0] add_67;
reg [39:0] add_68;
reg [39:0] add_69;
reg [39:0] add_70;
reg [39:0] add_71;
reg [39:0] add_72;
reg [39:0] add_73;
reg [39:0] add_74;
reg [39:0] add_75;
reg [39:0] add_76;
reg [39:0] add_77;
reg [39:0] add_78;
reg [39:0] add_79;

Delay_20bit d0(
	clk,
	in,
	z0
);

Delay_20bit d1(
  clk,
  z0,
  z1
);

Delay_20bit d2(
  clk,
  z1,
  z2
);

Delay_20bit d3(
  clk,
  z2,
  z3
);

Delay_20bit d4(
  clk,
  z3,
  z4
);

Delay_20bit d5(
  clk,
  z4,
  z5
);

Delay_20bit d6(
  clk,
  z5,
  z6
);

Delay_20bit d7(
  clk,
  z6,
  z7
);

Delay_20bit d8(
  clk,
  z7,
  z8
);

Delay_20bit d9(
  clk,
  z8,
  z9
);

Delay_20bit d10(
  clk,
  z9,
  z10
);

Delay_20bit d11(
  clk,
  z10,
  z11
);

Delay_20bit d12(
  clk,
  z11,
  z12
);

Delay_20bit d13(
  clk,
  z12,
  z13
);

Delay_20bit d14(
  clk,
  z13,
  z14
);

Delay_20bit d15(
  clk,
  z14,
  z15
);

Delay_20bit d16(
  clk,
  z15,
  z16
);

Delay_20bit d17(
  clk,
  z16,
  z17
);

Delay_20bit d18(
  clk,
  z17,
  z18
);

Delay_20bit d19(
  clk,
  z18,
  z19
);

Delay_20bit d20(
  clk,
  z19,
  z20
);

Delay_20bit d21(
  clk,
  z20,
  z21
);

Delay_20bit d22(
  clk,
  z21,
  z22
);

Delay_20bit d23(
  clk,
  z22,
  z23
);

Delay_20bit d24(
  clk,
  z23,
  z24
);

Delay_20bit d25(
  clk,
  z24,
  z25
);

Delay_20bit d26(
  clk,
  z25,
  z26
);

Delay_20bit d27(
  clk,
  z26,
  z27
);

Delay_20bit d28(
  clk,
  z27,
  z28
);

Delay_20bit d29(
  clk,
  z28,
  z29
);

Delay_20bit d30(
  clk,
  z29,
  z30
);

Delay_20bit d31(
  clk,
  z30,
  z31
);

Delay_20bit d32(
  clk,
  z31,
  z32
);

Delay_20bit d33(
  clk,
  z32,
  z33
);

Delay_20bit d34(
  clk,
  z33,
  z34
);

Delay_20bit d35(
  clk,
  z34,
  z35
);

Delay_20bit d36(
  clk,
  z35,
  z36
);

Delay_20bit d37(
  clk,
  z36,
  z37
);

Delay_20bit d38(
  clk,
  z37,
  z38
);

Delay_20bit d39(
  clk,
  z38,
  z39
);

Delay_20bit d40(
  clk,
  z39,
  z40
);

Delay_20bit d41(
  clk,
  z40,
  z41
);

Delay_20bit d42(
  clk,
  z41,
  z42
);

Delay_20bit d43(
  clk,
  z42,
  z43
);

Delay_20bit d44(
  clk,
  z43,
  z44
);

Delay_20bit d45(
  clk,
  z44,
  z45
);

Delay_20bit d46(
  clk,
  z45,
  z46
);

Delay_20bit d47(
  clk,
  z46,
  z47
);

Delay_20bit d48(
  clk,
  z47,
  z48
);

Delay_20bit d49(
  clk,
  z48,
  z49
);

Delay_20bit d50(
  clk,
  z49,
  z50
);

Delay_20bit d51(
  clk,
  z50,
  z51
);

Delay_20bit d52(
  clk,
  z51,
  z52
);

Delay_20bit d53(
  clk,
  z52,
  z53
);

Delay_20bit d54(
  clk,
  z53,
  z54
);

Delay_20bit d55(
  clk,
  z54,
  z55
);

Delay_20bit d56(
  clk,
  z55,
  z56
);

Delay_20bit d57(
  clk,
  z56,
  z57
);

Delay_20bit d58(
  clk,
  z57,
  z58
);

Delay_20bit d59(
  clk,
  z58,
  z59
);

Delay_20bit d60(
  clk,
  z59,
  z60
);

Delay_20bit d61(
  clk,
  z60,
  z61
);

Delay_20bit d62(
  clk,
  z61,
  z62
);

Delay_20bit d63(
  clk,
  z62,
  z63
);

Delay_20bit d64(
  clk,
  z63,
  z64
);

Delay_20bit d65(
  clk,
  z64,
  z65
);

Delay_20bit d66(
  clk,
  z65,
  z66
);

Delay_20bit d67(
  clk,
  z66,
  z67
);

Delay_20bit d68(
  clk,
  z67,
  z68
);

Delay_20bit d69(
  clk,
  z68,
  z69
);

Delay_20bit d70(
  clk,
  z69,
  z70
);

Delay_20bit d71(
  clk,
  z70,
  z71
);

Delay_20bit d72(
  clk,
  z71,
  z72
);

Delay_20bit d73(
  clk,
  z72,
  z73
);

Delay_20bit d74(
  clk,
  z73,
  z74
);

Delay_20bit d75(
  clk,
  z74,
  z75
);

Delay_20bit d76(
  clk,
  z75,
  z76
);

Delay_20bit d77(
  clk,
  z76,
  z77
);

Delay_20bit d78(
  clk,
  z77,
  z78
);

Delay_20bit d79(
  clk,
  z78,
  z79
);

Delay_20bit d80(
  clk,
  z79,
  z80
);

Delay_20bit d81(
  clk,
  z80,
  z81
);

Delay_20bit d82(
  clk,
  z81,
  z82
);

Delay_20bit d83(
  clk,
  z82,
  z83
);

Delay_20bit d84(
  clk,
  z83,
  z84
);

Delay_20bit d85(
  clk,
  z84,
  z85
);

Delay_20bit d86(
  clk,
  z85,
  z86
);

Delay_20bit d87(
  clk,
  z86,
  z87
);

Delay_20bit d88(
  clk,
  z87,
  z88
);

Delay_20bit d89(
  clk,
  z88,
  z89
);

Delay_20bit d90(
  clk,
  z89,
  z90
);

Delay_20bit d91(
  clk,
  z90,
  z91
);

Delay_20bit d92(
  clk,
  z91,
  z92
);

Delay_20bit d93(
  clk,
  z92,
  z93
);

Delay_20bit d94(
  clk,
  z93,
  z94
);

Delay_20bit d95(
  clk,
  z94,
  z95
);

Delay_20bit d96(
  clk,
  z95,
  z96
);

Delay_20bit d97(
  clk,
  z96,
  z97
);

Delay_20bit d98(
  clk,
  z97,
  z98
);

Delay_20bit d99(
  clk,
  z98,
  z99
);

Delay_20bit d100(
  clk,
  z99,
  z100
);

Delay_20bit d101(
  clk,
  z100,
  z101
);

Delay_20bit d102(
  clk,
  z101,
  z102
);

Delay_20bit d103(
  clk,
  z102,
  z103
);

Delay_20bit d104(
  clk,
  z103,
  z104
);

Delay_20bit d105(
  clk,
  z104,
  z105
);

Delay_20bit d106(
  clk,
  z105,
  z106
);

Delay_20bit d107(
  clk,
  z106,
  z107
);

Delay_20bit d108(
  clk,
  z107,
  z108
);

Delay_20bit d109(
  clk,
  z108,
  z109
);

Delay_20bit d110(
  clk,
  z109,
  z110
);

Delay_20bit d111(
  clk,
  z110,
  z111
);

Delay_20bit d112(
  clk,
  z111,
  z112
);

Delay_20bit d113(
  clk,
  z112,
  z113
);

Delay_20bit d114(
  clk,
  z113,
  z114
);

Delay_20bit d115(
  clk,
  z114,
  z115
);

Delay_20bit d116(
  clk,
  z115,
  z116
);

Delay_20bit d117(
  clk,
  z116,
  z117
);

Delay_20bit d118(
  clk,
  z117,
  z118
);

Delay_20bit d119(
  clk,
  z118,
  z119
);

Delay_20bit d120(
  clk,
  z119,
  z120
);

Delay_20bit d121(
  clk,
  z120,
  z121
);

Delay_20bit d122(
  clk,
  z121,
  z122
);

Delay_20bit d123(
  clk,
  z122,
  z123
);

Delay_20bit d124(
  clk,
  z123,
  z124
);

Delay_20bit d125(
  clk,
  z124,
  z125
);

Delay_20bit d126(
  clk,
  z125,
  z126
);

Delay_20bit d127(
  clk,
  z126,
  z127
);

Delay_20bit d128(
  clk,
  z127,
  z128
);

Delay_20bit d129(
  clk,
  z128,
  z129
);

Delay_20bit d130(
  clk,
  z129,
  z130
);

Delay_20bit d131(
  clk,
  z130,
  z131
);

Delay_20bit d132(
  clk,
  z131,
  z132
);

Delay_20bit d133(
  clk,
  z132,
  z133
);

Delay_20bit d134(
  clk,
  z133,
  z134
);

Delay_20bit d135(
  clk,
  z134,
  z135
);

Delay_20bit d136(
  clk,
  z135,
  z136
);

Delay_20bit d137(
  clk,
  z136,
  z137
);

Delay_20bit d138(
  clk,
  z137,
  z138
);

Delay_20bit d139(
  clk,
  z138,
  z139
);

Delay_20bit d140(
  clk,
  z139,
  z140
);

Delay_20bit d141(
  clk,
  z140,
  z141
);

Delay_20bit d142(
  clk,
  z141,
  z142
);

Delay_20bit d143(
  clk,
  z142,
  z143
);

Delay_20bit d144(
  clk,
  z143,
  z144
);

Delay_20bit d145(
  clk,
  z144,
  z145
);

Delay_20bit d146(
  clk,
  z145,
  z146
);

Delay_20bit d147(
  clk,
  z146,
  z147
);

Delay_20bit d148(
  clk,
  z147,
  z148
);

Delay_20bit d149(
  clk,
  z148,
  z149
);

Delay_20bit d150(
  clk,
  z149,
  z150
);

Delay_20bit d151(
  clk,
  z150,
  z151
);

Delay_20bit d152(
  clk,
  z151,
  z152
);

Delay_20bit d153(
  clk,
  z152,
  z153
);

Delay_20bit d154(
  clk,
  z153,
  z154
);

Delay_20bit d155(
  clk,
  z154,
  z155
);

Delay_20bit d156(
  clk,
  z155,
  z156
);

Delay_20bit d157(
  clk,
  z156,
  z157
);

Delay_20bit d158(
  clk,
  z157,
  z158
);

Delay_20bit d159(
  clk,
  z158,
  z159
);

Delay_20bit d160(
  clk,
  z159,
  z160
);

always @ (*) begin
	add0 <= z0 + z160;
	add1 <= z1 + z159;
	add2 <= z2 + z158;
	add3 <= z3 + z157;
	add4 <= z4 + z156;
	add5 <= z5 + z155;
	add6 <= z6 + z154;
	add7 <= z7 + z153;
	add8 <= z8 + z152;
	add9 <= z9 + z151;
	add10 <= z10 + z150;
	add11 <= z11 + z149;
	add12 <= z12 + z148;
	add13 <= z13 + z147;
	add14 <= z14 + z146;
	add15 <= z15 + z145;
	add16 <= z16 + z144;
	add17 <= z17 + z143;
	add18 <= z18 + z142;
	add19 <= z19 + z141;
	add20 <= z20 + z140;
	add21 <= z21 + z139;
	add22 <= z22 + z138;
	add23 <= z23 + z137;
	add24 <= z24 + z136;
	add25 <= z25 + z135;
	add26 <= z26 + z134;
	add27 <= z27 + z133;
	add28 <= z28 + z132;
	add29 <= z29 + z131;
	add30 <= z30 + z130;
	add31 <= z31 + z129;
	add32 <= z32 + z128;
	add33 <= z33 + z127;
	add34 <= z34 + z126;
	add35 <= z35 + z125;
	add36 <= z36 + z124;
	add37 <= z37 + z123;
	add38 <= z38 + z122;
	add39 <= z39 + z121;
	add40 <= z40 + z120;
	add41 <= z41 + z119;
	add42 <= z42 + z118;
	add43 <= z43 + z117;
	add44 <= z44 + z116;
	add45 <= z45 + z115;
	add46 <= z46 + z114;
	add47 <= z47 + z113;
	add48 <= z48 + z112;
	add49 <= z49 + z111;
	add50 <= z50 + z110;
	add51 <= z51 + z109;
	add52 <= z52 + z108;
	add53 <= z53 + z107;
	add54 <= z54 + z106;
	add55 <= z55 + z105;
	add56 <= z56 + z104;
	add57 <= z57 + z103;
	add58 <= z58 + z102;
	add59 <= z59 + z101;
	add60 <= z60 + z100;
	add61 <= z61 + z99;
	add62 <= z62 + z98;
	add63 <= z63 + z97;
	add64 <= z64 + z96;
	add65 <= z65 + z95;
	add66 <= z66 + z94;
	add67 <= z67 + z93;
	add68 <= z68 + z92;
	add69 <= z69 + z91;
	add70 <= z70 + z90;
	add71 <= z71 + z89;
	add72 <= z72 + z88;
	add73 <= z73 + z87;
	add74 <= z74 + z86;
	add75 <= z75 + z85;
	add76 <= z76 + z84;
	add77 <= z77 + z83;
	add78 <= z78 + z82;
	add79 <= z79 + z81;
	
	mult0 <= add0 * h0;
	mult1 <= add1 * h1;
	mult2 <= add2 * h2;
	mult3 <= add3 * h3;
	mult4 <= add4 * h4;
	mult5 <= add5 * h5;
	mult6 <= add6 * h6;
	mult7 <= add7 * h7;
	mult8 <= add8 * h8;
	mult9 <= add9 * h9;
	mult10 <= add10 * h10;
	mult11 <= add11 * h11;
	mult12 <= add12 * h12;
	mult13 <= add13 * h13;
	mult14 <= add14 * h14;
	mult15 <= add15 * h15;
	mult16 <= add16 * h16;
	mult17 <= add17 * h17;
	mult18 <= add18 * h18;
	mult19 <= add19 * h19;
	mult20 <= add20 * h20;
	mult21 <= add21 * h21;
	mult22 <= add22 * h22;
	mult23 <= add23 * h23;
	mult24 <= add24 * h24;
	mult25 <= add25 * h25;
	mult26 <= add26 * h26;
	mult27 <= add27 * h27;
	mult28 <= add28 * h28;
	mult29 <= add29 * h29;
	mult30 <= add30 * h30;
	mult31 <= add31 * h31;
	mult32 <= add32 * h32;
	mult33 <= add33 * h33;
	mult34 <= add34 * h34;
	mult35 <= add35 * h35;
	mult36 <= add36 * h36;
	mult37 <= add37 * h37;
	mult38 <= add38 * h38;
	mult39 <= add39 * h39;
	mult40 <= add40 * h40;
	mult41 <= add41 * h41;
	mult42 <= add42 * h42;
	mult43 <= add43 * h43;
	mult44 <= add44 * h44;
	mult45 <= add45 * h45;
	mult46 <= add46 * h46;
	mult47 <= add47 * h47;
	mult48 <= add48 * h48;
	mult49 <= add49 * h49;
	mult50 <= add50 * h50;
	mult51 <= add51 * h51;
	mult52 <= add52 * h52;
	mult53 <= add53 * h53;
	mult54 <= add54 * h54;
	mult55 <= add55 * h55;
	mult56 <= add56 * h56;
	mult57 <= add57 * h57;
	mult58 <= add58 * h58;
	mult59 <= add59 * h59;
	mult60 <= add60 * h60;
	mult61 <= add61 * h61;
	mult62 <= add62 * h62;
	mult63 <= add63 * h63;
	mult64 <= add64 * h64;
	mult65 <= add65 * h65;
	mult66 <= add66 * h66;
	mult67 <= add67 * h67;
	mult68 <= add68 * h68;
	mult69 <= add69 * h69;
	mult70 <= add70 * h70;
	mult71 <= add71 * h71;
	mult72 <= add72 * h72;
	mult73 <= add73 * h73;
	mult74 <= add74 * h74;
	mult75 <= add75 * h75;
	mult76 <= add76 * h76;
	mult77 <= add77 * h77;
	mult78 <= add78 * h78;
	mult79 <= add79 * h79;
	mult80 <= z80 * h80;
	
	add_0 <= mult80 + mult79;
	add_1 <= add_0 + mult78;
	add_2 <= add_1 + mult77;
	add_3 <= add_2 + mult76;
	add_4 <= add_3 + mult75;
	add_5 <= add_4 + mult74;
	add_6 <= add_5 + mult73;
	add_7 <= add_6 + mult72;
	add_8 <= add_7 + mult71;
	add_9 <= add_8 + mult70;
	add_10 <= add_9 + mult69;
	add_11 <= add_10 + mult68;
	add_12 <= add_11 + mult67;
	add_13 <= add_12 + mult66;
	add_14 <= add_13 + mult65;
	add_15 <= add_14 + mult64;
	add_16 <= add_15 + mult63;
	add_17 <= add_16 + mult62;
	add_18 <= add_17 + mult61;
	add_19 <= add_18 + mult60;
	add_20 <= add_19 + mult59;
	add_21 <= add_20 + mult58;
	add_22 <= add_21 + mult57;
	add_23 <= add_22 + mult56;
	add_24 <= add_23 + mult55;
	add_25 <= add_24 + mult54;
	add_26 <= add_25 + mult53;
	add_27 <= add_26 + mult52;
	add_28 <= add_27 + mult51;
	add_29 <= add_28 + mult50;
	add_30 <= add_29 + mult49;
	add_31 <= add_30 + mult48;
	add_32 <= add_31 + mult47;
	add_33 <= add_32 + mult46;
	add_34 <= add_33 + mult45;
	add_35 <= add_34 + mult44;
	add_36 <= add_35 + mult43;
	add_37 <= add_36 + mult42;
	add_38 <= add_37 + mult41;
	add_39 <= add_38 + mult40;
	add_40 <= add_39 + mult39;
	add_41 <= add_40 + mult38;
	add_42 <= add_41 + mult37;
	add_43 <= add_42 + mult36;
	add_44 <= add_43 + mult35;
	add_45 <= add_44 + mult34;
	add_46 <= add_45 + mult33;
	add_47 <= add_46 + mult32;
	add_48 <= add_47 + mult31;
	add_49 <= add_48 + mult30;
	add_50 <= add_49 + mult29;
	add_51 <= add_50 + mult28;
	add_52 <= add_51 + mult27;
	add_53 <= add_52 + mult26;
	add_54 <= add_53 + mult25;
	add_55 <= add_54 + mult24;
	add_56 <= add_55 + mult23;
	add_57 <= add_56 + mult22;
	add_58 <= add_57 + mult21;
	add_59 <= add_58 + mult20;
	add_60 <= add_59 + mult19;
	add_61 <= add_60 + mult18;
	add_62 <= add_61 + mult17;
	add_63 <= add_62 + mult16;
	add_64 <= add_63 + mult15;
	add_65 <= add_64 + mult14;
	add_66 <= add_65 + mult13;
	add_67 <= add_66 + mult12;
	add_68 <= add_67 + mult11;
	add_69 <= add_68 + mult10;
	add_70 <= add_69 + mult9;
	add_71 <= add_70 + mult8;
	add_72 <= add_71 + mult7;
	add_73 <= add_72 + mult6;
	add_74 <= add_73 + mult5;
	add_75 <= add_74 + mult4;
	add_76 <= add_75 + mult3;
	add_77 <= add_76 + mult2;
	add_78 <= add_77 + mult1;
	add_79 <= add_78 + mult0;
end

assign out = add_79;

endmodule