module mux2bitS(
	input Sel,
	input In1,
	input In2,
	
	output Out

);

always @(Sel) begin


end



endmodule
