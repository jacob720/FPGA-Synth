module DE2_load_program( A, B, Out );

input A;
input B;

output Out;

and(Out, A, B);

endmodule
